/*
CPEN311 Lab 2: Circles and Triangles
Ansh Madaan (8399574) & Rishi Upath (18259374)
October 27, 2025

SYN Testbench for task4 Module
Purpose: Tests task4 modules output signals by implementing a reference reuleaux triangle algorithm and comparing.
         Checks for vga_x, vga_y, vga_plot, and colour.
*/

`timescale 1ps/1ps

module tb_syn_task4();

    reg tb_CLOCK_50;
    reg [3:0] tb_KEY;
    reg [9:0] tb_SW; 
    wire [9:0] tb_LEDR;
    wire [6:0] tb_HEX0, tb_HEX1, tb_HEX2, tb_HEX3, tb_HEX4, tb_HEX5;
    wire [7:0] tb_VGA_R, tb_VGA_G, tb_VGA_B, tb_VGA_X;
    wire [6:0] tb_VGA_Y;
    wire [2:0] tb_VGA_COLOUR;
    wire tb_VGA_HS, tb_VGA_VS, tb_VGA_CLK, tb_VGA_PLOT;
    
    reg err;
    
    //instantiate task4 module
    task4 DUT(.CLOCK_50(tb_CLOCK_50), .KEY(tb_KEY), .SW(tb_SW), .LEDR(tb_LEDR), .HEX0(tb_HEX0),
             .HEX1(tb_HEX1), .HEX2(tb_HEX2), .HEX3(tb_HEX3), .HEX4(tb_HEX4), .HEX5(tb_HEX5),
             .VGA_R(tb_VGA_R), .VGA_G(tb_VGA_G), .VGA_B(tb_VGA_B),
             .VGA_HS(tb_VGA_HS), .VGA_VS(tb_VGA_VS), .VGA_CLK(tb_VGA_CLK),
             .VGA_X(tb_VGA_X), .VGA_Y(tb_VGA_Y),
             .VGA_COLOUR(tb_VGA_COLOUR), .VGA_PLOT(tb_VGA_PLOT));

    //local regs to compute pixels positions to draw
    reg signed [7:0] expected_offset_y;
    reg signed [7:0] expected_offset_x;
    reg signed [8:0] expected_crit;

    reg signed [8:0] signed_centre_x, expected_vga_x;
    reg signed [8:0] signed_centre_y, expected_vga_y;
    reg [7:0] tb_diameter;

    real expected_top_centre_x, expected_left_centre_x, expected_right_centre_x;
    real expected_top_centre_y, expected_left_centre_y, expected_right_centre_y;

    reg expected_vga_plot;

    //signed version of centre x and y
    assign signed_centre_x = 9'sd80;
    assign signed_centre_y = 9'sd60;

    //diameter
    assign tb_diameter = 8'd80;

    //task checker for fillscreen module, checks x and y position, colour, and plot
    task fillscreen_checker;
        
        input [7:0] x_expected;
        input [6:0] y_expected;
        input [2:0] colour_expected;
        input vga_plot_expected;

        begin
            
            if (tb_syn_task4.DUT.VGA_X != x_expected) begin
                $display("ERROR, x position is %b, expected %b", tb_syn_task4.DUT.VGA_X, x_expected);
                err = 1'b1;
            end
            if (tb_syn_task4.DUT.VGA_Y != y_expected) begin
                $display("ERROR, y position is %b, expected %b", tb_syn_task4.DUT.VGA_Y, y_expected);
                err = 1'b1;
            end
            if (tb_syn_task4.DUT.VGA_COLOUR != colour_expected) begin
                $display("ERROR, colour is %b, expected %b", tb_syn_task4.DUT.VGA_COLOUR, colour_expected);
                err = 1'b1;
            end
            if (tb_syn_task4.DUT.VGA_PLOT != vga_plot_expected) begin
                $display("ERROR, vga_plot is %b, expected %b", tb_syn_task4.DUT.VGA_PLOT, vga_plot_expected);
                err = 1'b1;
            end

        end
    endtask
    
    //task checker for drawing circle, tests vga_x, vga_y, vga_plot, crit, offsets, start, and done signals
    task reuleaux_checker;

        begin
            //initialize local parameters
            expected_offset_y = 7'd0;
            expected_offset_x = tb_diameter;
            expected_crit = 9'sd1 - $signed(tb_diameter);

            //compute expected centres 
            expected_top_centre_x = signed_centre_x;
            expected_top_centre_y = signed_centre_y - tb_diameter * ($sqrt(3.0)/3.0);
            expected_left_centre_x = signed_centre_x - tb_diameter / 2;
            expected_left_centre_y = signed_centre_y + tb_diameter * ($sqrt(3.0)/6.0);
            expected_right_centre_x = signed_centre_x + tb_diameter / 2;
            expected_right_centre_y = signed_centre_y + tb_diameter * ($sqrt(3.0)/6.0);

            while (expected_offset_y <= expected_offset_x) begin 

                @(posedge tb_CLOCK_50); #1;
                //octant 8 test
                expected_vga_x = int'(expected_left_centre_x) + expected_offset_x;
                expected_vga_y = int'(expected_left_centre_y) - expected_offset_y; #1;
                
                //checking vga_x
                $display("Checking vga_x, octant 8");
                if (tb_syn_task4.DUT.VGA_X != expected_vga_x[7:0]) begin 
                    err = 1'b1;
                    $display("vga_x is %b, expected vga_x is %b", tb_syn_task4.DUT.VGA_X, expected_vga_x);
                end

                //checking vga_y
                $display("Checking vga_y, octant 8");
                if (tb_syn_task4.DUT.VGA_Y != expected_vga_y[6:0]) begin
                    err = 1'b1;
                    $display("vga_y is %b, expected vga_y is %b", tb_syn_task4.DUT.VGA_Y, expected_vga_y);
                end

                //determine expected plot depending on boundary condition
                if (expected_vga_x < 9'sd0 || expected_vga_x > 9'sd159)
                    expected_vga_plot = 1'b0;
                else if (expected_vga_y < 9'sd0 || expected_vga_y > 9'sd119)
                    expected_vga_plot = 1'b0;
                else if ((expected_vga_x > int'(expected_right_centre_x)) || (expected_vga_x < int'(expected_top_centre_x)) || (expected_vga_y < int'(expected_top_centre_y)) || (expected_vga_y > int'(expected_right_centre_y))) 
                    expected_vga_plot = 1'b0;
                else 
                    expected_vga_plot = 1'b1;

                //check if plot is high
                $display("Checking plot signal");
                if (tb_syn_task4.DUT.VGA_PLOT != expected_vga_plot) begin
                    err = 1'b1;
                    $display("vga_plot is %b, expected %b",tb_syn_task4.DUT.VGA_PLOT, expected_vga_plot);
                end



                @(posedge tb_CLOCK_50); #1;
                //octant 7 test
                expected_vga_x = int'(expected_left_centre_x) + expected_offset_y;
                expected_vga_y = int'(expected_left_centre_y) - expected_offset_x; #1;
                
                $display("Checking vga_x, octant 7");
                if (tb_syn_task4.DUT.VGA_X != expected_vga_x[7:0]) begin 
                    err = 1'b1;
                    $display("vga_x is %b, expected vga_x is %b", tb_syn_task4.DUT.VGA_X, expected_vga_x);
                end

                $display("Checking vga_y, octant 7");
                if (tb_syn_task4.DUT.VGA_Y != expected_vga_y[6:0]) begin
                    err = 1'b1;
                    $display("vga_y is %b, expected vga_y is %b", tb_syn_task4.DUT.VGA_Y, expected_vga_y);
                end

                //determine expected plot depending on boundary condition
                if (expected_vga_x < 9'sd0 || expected_vga_x > 9'sd159)
                    expected_vga_plot = 1'b0;
                else if (expected_vga_y < 9'sd0 || expected_vga_y > 9'sd119)
                    expected_vga_plot = 1'b0;
                else if ((expected_vga_x > int'(expected_right_centre_x)) || (expected_vga_x < int'(expected_top_centre_x)) || (expected_vga_y < int'(expected_top_centre_y)) || (expected_vga_y > int'(expected_right_centre_y))) 
                    expected_vga_plot = 1'b0;
                else 
                    expected_vga_plot = 1'b1;

                //check if plot is high
                $display("Checking plot signal");
                if (tb_syn_task4.DUT.VGA_PLOT != expected_vga_plot) begin
                    err = 1'b1;
                    $display("vga_plot is %b, expected %b",tb_syn_task4.DUT.VGA_PLOT, expected_vga_plot);
                end



                @(posedge tb_CLOCK_50); #1;
                //octant 6 test
                expected_vga_x = int'(expected_right_centre_x) - expected_offset_y;
                expected_vga_y = int'(expected_right_centre_y) - expected_offset_x; #1;
                
                $display("Checking vga_x, octant 6");
                if (tb_syn_task4.DUT.VGA_X != expected_vga_x[7:0]) begin 
                    err = 1'b1;
                    $display("vga_x is %b, expected vga_x is %b", tb_syn_task4.DUT.VGA_X, expected_vga_x);
                end

                $display("Checking vga_y, octant 6");
                if (tb_syn_task4.DUT.VGA_Y != expected_vga_y[6:0]) begin
                    err = 1'b1;
                    $display("vga_y is %b, expected vga_y is %b", tb_syn_task4.DUT.VGA_Y, expected_vga_y);
                end

                //determine expected plot depending on boundary condition
                if (expected_vga_x < 9'sd0 || expected_vga_x > 9'sd159)
                    expected_vga_plot = 1'b0;
                else if (expected_vga_y < 9'sd0 || expected_vga_y > 9'sd119)
                    expected_vga_plot = 1'b0;
                else if ((expected_vga_x > int'(expected_top_centre_x)) || (expected_vga_x < int'(expected_left_centre_x)) || (expected_vga_y < int'(expected_top_centre_y)) || (expected_vga_y > int'(expected_left_centre_y))) 
                    expected_vga_plot = 1'b0;
                else 
                    expected_vga_plot = 1'b1;

                //check if plot is high
                $display("Checking plot signal");
                if (tb_syn_task4.DUT.VGA_PLOT != expected_vga_plot) begin
                    err = 1'b1;
                    $display("vga_plot is %b, expected %b",tb_syn_task4.DUT.VGA_PLOT, expected_vga_plot);
                end



                @(posedge tb_CLOCK_50); #1;
                //octant 5 test
                expected_vga_x = int'(expected_right_centre_x) - expected_offset_x;
                expected_vga_y = int'(expected_right_centre_y) - expected_offset_y; #1;
                
                $display("Checking vga_x, octant 5");
                if (tb_syn_task4.DUT.VGA_X != expected_vga_x[7:0]) begin 
                    err = 1'b1;
                    $display("vga_x is %b, expected vga_x is %b", tb_syn_task4.DUT.VGA_X, expected_vga_x);
                end

                $display("Checking vga_y, octant 5");
                if (tb_syn_task4.DUT.VGA_Y != expected_vga_y[6:0]) begin
                    err = 1'b1;
                    $display("vga_y is %b, expected vga_y is %b", tb_syn_task4.DUT.VGA_Y, expected_vga_y);
                end

                //determine expected plot depending on boundary condition
                if (expected_vga_x < 9'sd0 || expected_vga_x > 9'sd159)
                    expected_vga_plot = 1'b0;
                else if (expected_vga_y < 9'sd0 || expected_vga_y > 9'sd119)
                    expected_vga_plot = 1'b0;
                else if ((expected_vga_x > int'(expected_top_centre_x)) || (expected_vga_x < int'(expected_left_centre_x)) || (expected_vga_y < int'(expected_top_centre_y)) || (expected_vga_y > int'(expected_left_centre_y))) 
                    expected_vga_plot = 1'b0;
                else 
                    expected_vga_plot = 1'b1;

                //check if plot is high
                $display("Checking plot signal");
                if (tb_syn_task4.DUT.VGA_PLOT != expected_vga_plot) begin
                    err = 1'b1;
                    $display("vga_plot is %b, expected %b",tb_syn_task4.DUT.VGA_PLOT, expected_vga_plot);
                end



                @(posedge tb_CLOCK_50); #1;
                //octant 3 test
                expected_vga_x = int'(expected_top_centre_x) - expected_offset_y;
                expected_vga_y = int'(expected_top_centre_y) + expected_offset_x; #1;

                $display("Checking vga_x, octant 3");
                if (tb_syn_task4.DUT.VGA_X != expected_vga_x[7:0]) begin 
                    err = 1'b1;
                    $display("vga_x is %b, expected vga_x is %b", tb_syn_task4.DUT.VGA_X, expected_vga_x);
                end

                $display("Checking vga_y, octant 3");
                if (tb_syn_task4.DUT.VGA_Y != expected_vga_y[6:0]) begin
                    err = 1'b1;
                    $display("vga_y is %b, expected vga_y is %b", tb_syn_task4.DUT.VGA_Y, expected_vga_y);
                end

                //determine expected plot depending on boundary condition
                if (expected_vga_x < 9'sd0 || expected_vga_x > 9'sd159)
                    expected_vga_plot = 1'b0;
                else if (expected_vga_y < 9'sd0 || expected_vga_y > 9'sd119)
                    expected_vga_plot = 1'b0;
                else if ((expected_vga_x > int'(expected_right_centre_x)) || (expected_vga_x < int'(expected_left_centre_x)) || (expected_vga_y < int'(expected_right_centre_y)))
                    expected_vga_plot = 1'b0;
                else 
                    expected_vga_plot = 1'b1;

                //check if plot is high
                $display("Checking plot signal");
                if (tb_syn_task4.DUT.VGA_PLOT != expected_vga_plot) begin
                    err = 1'b1;
                    $display("vga_plot is %b, expected %b",tb_syn_task4.DUT.VGA_PLOT, expected_vga_plot);
                end



                @(posedge tb_CLOCK_50); #1;
                //octant 2 test
                expected_vga_x = int'(expected_top_centre_x) + expected_offset_y;
                expected_vga_y = int'(expected_top_centre_y) + expected_offset_x; #1;
                
                $display("Checking vga_x, octant 2");
                if (tb_syn_task4.DUT.VGA_X != expected_vga_x[7:0]) begin 
                    err = 1'b1;
                    $display("vga_x is %b, expected vga_x is %b", tb_syn_task4.DUT.VGA_X, expected_vga_x);
                end

                $display("Checking vga_y, octant 2");
                if (tb_syn_task4.DUT.VGA_Y != expected_vga_y[6:0]) begin
                    err = 1'b1;
                    $display("vga_y is %b, expected vga_y is %b", tb_syn_task4.DUT.VGA_Y, expected_vga_y);
                end  

                //determine expected plot depending on boundary condition
                if (expected_vga_x < 9'sd0 || expected_vga_x > 9'sd159)
                    expected_vga_plot = 1'b0;
                else if (expected_vga_y < 9'sd0 || expected_vga_y > 9'sd119)
                    expected_vga_plot = 1'b0;
                else if ((expected_vga_x > int'(expected_right_centre_x)) || (expected_vga_x < int'(expected_left_centre_x)) || (expected_vga_y < int'(expected_right_centre_y)))
                    expected_vga_plot = 1'b0;
                else 
                    expected_vga_plot = 1'b1;

                //check if plot is high
                $display("Checking plot signal");
                if (tb_syn_task4.DUT.VGA_PLOT != expected_vga_plot) begin
                    err = 1'b1;
                    $display("vga_plot is %b, expected %b",tb_syn_task4.DUT.VGA_PLOT, expected_vga_plot);
                end

                //changing offset_y, offset_x, and crit according to reuleauxdrawing algorithm 
                expected_offset_y = expected_offset_y + 8'sd1;

                if (expected_crit <= 9'sd0)
                    expected_crit = expected_crit + 9'sd2 * $signed(expected_offset_y) + 9'sd1;
                else begin
                    expected_offset_x = expected_offset_x - 8'sd1;
                    expected_crit = expected_crit + 9'sd2 * ($signed(expected_offset_y) - $signed(expected_offset_x)) + 9'sd1;
                end

            end
            
            @(posedge tb_CLOCK_50); #1;
            @(posedge tb_CLOCK_50); #1;

            //check if plot is low
            $display("Checking plot signal");
            if (tb_syn_task4.DUT.VGA_PLOT != 1'b0) begin
            err = 1'b1;
            $display("vga_plot is %b, expected 0",tb_syn_task4.DUT.VGA_PLOT);
            end
            
        end

    endtask 

    //initializing tb_CLOCK_50 for each pixel
    initial begin 
        tb_CLOCK_50 = 1'b0; #10; 

        forever begin
            tb_CLOCK_50 = 1'b1; #10;
            tb_CLOCK_50 = 1'b0; #10;
        end
    end

    //block to test fillscreen and circle together
    initial begin
        err = 1'b0;

        //assert reset
        tb_KEY[3] = 1'b0; #20;
        tb_KEY[3] = 1'b1; #5;

        @(posedge tb_CLOCK_50); #1;

        //fillscreen colours the entire screen black

        //check colour
        $display("Checking colour is black");
        if (tb_syn_task4.DUT.VGA_COLOUR != 3'b000) begin 
            err = 1'b1;
            $display("colour is %b, expected 000 (black)", tb_syn_task4.DUT.VGA_COLOUR);
        end

        //check position and colour of every pixel as well as correct plot signal
        for (integer i = 0; i <= 159; i++) begin
            for (integer j = 0; j <= 119; j++) begin 
                //account for extra increment of y after reset
                if (i == 0 && j == 0) 
                    j++;

                $display("Start time is, %0t", $time);
                fillscreen_checker(i, j, 3'b000, 1'b1);
                #20;
            end 
        end

        //check for fillscreen_start, reuleaux_start
        @(posedge tb_CLOCK_50); #1;

        //check colour
        $display("Checking colour is green");
        if (tb_syn_task4.DUT.VGA_COLOUR != 3'b010) begin 
            err = 1'b1;
            $display("colour is %b, expected 010 (green)", tb_syn_task4.DUT.VGA_COLOUR);
        end

        //checking reuleaux
        $display("Testing reuleaux with radius: 80, centre: (80,60) at: %0t", $time);
        reuleaux_checker();

        //display error or passed message 
        if(err)
            $display("Some cases FAILED :(");
        else 
            $display("All cases PASSED :)");
            
        $stop;

    end

endmodule: tb_syn_task4
